module float_adder(
    input           clk,
    input   [31:0]  a,
    output  [31:0]  b);

    reg     

endmodule